library verilog;
use verilog.vl_types.all;
entity LATCH_SR_NOR_vlg_vec_tst is
end LATCH_SR_NOR_vlg_vec_tst;
