library verilog;
use verilog.vl_types.all;
entity Practica_2_vlg_sample_tst is
    port(
        C               : in     vl_logic;
        E               : in     vl_logic;
        S               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Practica_2_vlg_sample_tst;
