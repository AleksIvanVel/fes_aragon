library verilog;
use verilog.vl_types.all;
entity LATCH_TIPO_NAND_vlg_sample_tst is
    port(
        Rn              : in     vl_logic;
        Sn              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end LATCH_TIPO_NAND_vlg_sample_tst;
