library verilog;
use verilog.vl_types.all;
entity SM_CONTADOR_vlg_vec_tst is
end SM_CONTADOR_vlg_vec_tst;
