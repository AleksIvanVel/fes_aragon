library verilog;
use verilog.vl_types.all;
entity Practica_2_vlg_check_tst is
    port(
        A               : in     vl_logic;
        R               : in     vl_logic;
        V               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Practica_2_vlg_check_tst;
