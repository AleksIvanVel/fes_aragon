library verilog;
use verilog.vl_types.all;
entity Practica_2_vlg_vec_tst is
end Practica_2_vlg_vec_tst;
