library verilog;
use verilog.vl_types.all;
entity CONTADOR_vlg_vec_tst is
end CONTADOR_vlg_vec_tst;
