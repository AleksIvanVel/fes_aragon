library verilog;
use verilog.vl_types.all;
entity Practica_2 is
    port(
        S               : in     vl_logic;
        E               : in     vl_logic;
        C               : in     vl_logic;
        R               : out    vl_logic;
        A               : out    vl_logic;
        V               : out    vl_logic
    );
end Practica_2;
