// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
// Created on Wed Mar 13 09:33:53 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module SM_CONTADOR (
    reset,clock,input1,
    output1,output2,output3);

    input reset;
    input clock;
    input input1;
    tri0 reset;
    tri0 input1;
    output output1;
    output output2;
    output output3;
    reg output1;
    reg output2;
    reg output3;
    reg [7:0] fstate;
    reg [7:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state8=4,state6=5,state7=6,state5=7;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or input1)
    begin
        if (reset) begin
            reg_fstate <= state1;
            output1 <= 1'b0;
            output2 <= 1'b0;
            output3 <= 1'b0;
        end
        else begin
            output1 <= 1'b0;
            output2 <= 1'b0;
            output3 <= 1'b0;
            case (fstate)
                state1: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state8;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    output2 <= 1'b0;

                    output3 <= 1'b0;

                    output1 <= 1'b0;
                end
                state2: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state1;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    output2 <= 1'b0;

                    output3 <= 1'b1;

                    output1 <= 1'b0;
                end
                state3: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state2;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    output2 <= 1'b1;

                    output3 <= 1'b0;

                    output1 <= 1'b0;
                end
                state4: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state3;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    output2 <= 1'b1;

                    output3 <= 1'b1;

                    output1 <= 1'b0;
                end
                state8: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state1;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state7;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state8;

                    output2 <= 1'b1;

                    output3 <= 1'b1;

                    output1 <= 1'b1;
                end
                state6: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state5;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state7;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state6;

                    output2 <= 1'b0;

                    output3 <= 1'b1;

                    output1 <= 1'b1;
                end
                state7: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state6;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state7;

                    output2 <= 1'b1;

                    output3 <= 1'b0;

                    output1 <= 1'b1;
                end
                state5: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state4;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    output2 <= 1'b0;

                    output3 <= 1'b0;

                    output1 <= 1'b1;
                end
                default: begin
                    output1 <= 1'bx;
                    output2 <= 1'bx;
                    output3 <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM_CONTADOR
