library verilog;
use verilog.vl_types.all;
entity LATCH_TIPO_D_vlg_vec_tst is
end LATCH_TIPO_D_vlg_vec_tst;
